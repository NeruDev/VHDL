---------------------------------------------------------------------
-- LIBRERIAS
---------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
--USE ieee.numeric_std.all;

---------------------------------------------------------------------
-- ENTIDAD
---------------------------------------------------------------------
ENTITY BASE IS

  PORT (
    A : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
    X : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END ENTITY BASE;

---------------------------------------------------------------------
-- ARQUITECTURA
---------------------------------------------------------------------
ARCHITECTURE UNO OF BASE IS

BEGIN

END ARCHITECTURE UNO;