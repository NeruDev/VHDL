---------------------------------------------------------------------
-- PLANTILLA REDUCIDA VHDL
---------------------------------------------------------------------

---------------------------------------------------------------------
-- LIBRERIAS
---------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
--USE ieee.numeric_std.all;

---------------------------------------------------------------------
-- ENTIDAD
---------------------------------------------------------------------
ENTITY plantilla_design_testbench IS
   GENERIC (
      G_DATA_WIDTH  : INTEGER := 8
   );
   PORT (
      i_data_a : IN  STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0);
      i_data_b : IN  STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0);
      i_sel    : IN  STD_LOGIC;
      o_data   : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0)
   );
END ENTITY plantilla_design_testbench;

---------------------------------------------------------------------
-- ARQUITECTURA
---------------------------------------------------------------------
ARCHITECTURE behavioral OF plantilla_design_testbench IS

   -------------------------------------------------------------------
   -- CONSTANTES
   -------------------------------------------------------------------

   -------------------------------------------------------------------
   -- SEÑALES
   -------------------------------------------------------------------

   -------------------------------------------------------------------
   -- COMPONENTES
   -------------------------------------------------------------------

   -------------------------------------------------------------------
   -- FUNCIONES Y PROCEDIMIENTOS
   -------------------------------------------------------------------

BEGIN

   -------------------------------------------------------------------
   -- ASIGNACIONES CONCURRENTES
   -------------------------------------------------------------------

   -------------------------------------------------------------------
   -- PROCESOS
   -------------------------------------------------------------------

END ARCHITECTURE behavioral;